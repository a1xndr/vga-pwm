WARNING:ProjectMgmt - File /home/alxndr/Develpoment/FPGA/vga_test/vga_vhdl.prj is missing.
